// `include "data_structures.sv"

// module extract_reg(
//     input logic [31:0] insnbits.
//     input logic [`OPCODE_SIZE-1:0] op,
//     output logic [`GPR_IDX_SIZE-1:0] src1,
//     output logic [`GPR_IDX_SIZE-1:0] src2,
//     output logic [`GPR_IDX_SIZE-1:0] dst,
// );

//     casez(op)
    

//     endcase

// endmodule